module rom	(
input		wire	[7:0]		addr,
output	reg	[26:0]	data
);

always @*
	case(addr)
		8'h00		:	data	=	27'b000000000000000001000000000; //FETCH
		8'h01		:	data	=	27'b000110001000000000000100000;
		8'h02		:	data	=	27'b000000000000000100001010000;
		8'h03		:	data	=	27'b000000000000000000000000000;
		8'h04		:	data	=	27'b000000000000000000000000000;
		8'h05		:	data	=	27'b000000000000000000000000000;
		8'h06		:	data	=	27'b000000000000000000000000000;
		8'h07		:	data	=	27'b000000000000000000000000000;
		8'h08		:	data	=	27'b001000001011111010000010000; //MOV ACC A
		8'h09		:	data	=	27'b000000000000000000000000000;
		8'h0A		:	data	=	27'b000000000000000000000000000;
		8'h0B		:	data	=	27'b000000000000000000000000000;
		8'h0C		:	data	=	27'b000000000000000000000000000;
		8'h0D		:	data	=	27'b000000000000000000000000000;
		8'h0E		:	data	=	27'b000000000000000000000000000;
		8'h0F		:	data	=	27'b000000000000000000000000000;
		8'h10		:	data	=	27'b001000001111011010000010000; //MOV A ACC
		8'h11		:	data	=	27'b000000000000000000000000000;
		8'h12		:	data	=	27'b000000000000000000000000000;
		8'h13		:	data	=	27'b000000000000000000000000000;
		8'h14		:	data	=	27'b000000000000000000000000000;
		8'h15		:	data	=	27'b000000000000000000000000000;
		8'h16		:	data	=	27'b000000000000000000000000000;
		8'h17		:	data	=	27'b000000000000000000000000000;
		8'h18		:	data	=	27'b000000000000000001000000000; //MOV ACC CTE
		8'h19		:	data	=	27'b000110001000000000000100000;
		8'h1A		:	data	=	27'b000000001000111010001010000;
		8'h1B		:	data	=	27'b000000000000000000000000000;
		8'h1C		:	data	=	27'b000000000000000000000000000;
		8'h1D		:	data	=	27'b000000000000000000000000000;
		8'h1E		:	data	=	27'b000000000000000000000000000;
		8'h1F		:	data	=	27'b000000000000000000000000000;
		8'h20		:	data	=	27'b000000000010000001000000000; //MOV ACC [DPTR]
		8'h21		:	data	=	27'b000000000000000000000100000;
		8'h22		:	data	=	27'b000000001000111010001010000;
		8'h23		:	data	=	27'b000000000000000000000000000;
		8'h24		:	data	=	27'b000000000000000000000000000;
		8'h25		:	data	=	27'b000000000000000000000000000;
		8'h26		:	data	=	27'b000000000000000000000000000;
		8'h27		:	data	=	27'b000000000000000000000000000;
		8'h28		:	data	=	27'b001000001111010010000010000; //MOV DPTR ACC
		8'h29		:	data	=	27'b000000000000000000000000000;
		8'h2A		:	data	=	27'b000000000000000000000000000;
		8'h2B		:	data	=	27'b000000000000000000000000000;
		8'h2C		:	data	=	27'b000000000000000000000000000;
		8'h2D		:	data	=	27'b000000000000000000000000000;
		8'h2E		:	data	=	27'b000000000000000000000000000;
		8'h2F		:	data	=	27'b000000000000000000000000000;
		8'h30		:	data	=	27'b000000000111000000000100000; //MOV [DPTR] ACC
		8'h31		:	data	=	27'b000000000010000001000000000;
		8'h32		:	data	=	27'b001000000000000010010010000;
		8'h33		:	data	=	27'b000000000000000000000000000;
		8'h34		:	data	=	27'b000000000000000000000000000;
		8'h35		:	data	=	27'b000000000000000000000000000;
		8'h36		:	data	=	27'b000000000000000000000000000;
		8'h37		:	data	=	27'b000000000000000000000000000;
		8'h38		:	data	=	27'b001001001111111010000010000; //INV ACC
		8'h39		:	data	=	27'b000000000000000000000000000;
		8'h3A		:	data	=	27'b000000000000000000000000000;
		8'h3B		:	data	=	27'b000000000000000000000000000;
		8'h3C		:	data	=	27'b000000000000000000000000000;
		8'h3D		:	data	=	27'b000000000000000000000000000;
		8'h3E		:	data	=	27'b000000000000000000000000000;
		8'h3F		:	data	=	27'b000000000000000000000000000;
		8'h40		:	data	=	27'b001010001011111010000010000; //AND ACC A
		8'h41		:	data	=	27'b000000000000000000000000000;
		8'h42		:	data	=	27'b000000000000000000000000000;
		8'h43		:	data	=	27'b000000000000000000000000000;
		8'h44		:	data	=	27'b000000000000000000000000000;
		8'h45		:	data	=	27'b000000000000000000000000000;
		8'h46		:	data	=	27'b000000000000000000000000000;
		8'h47		:	data	=	27'b000000000000000000000000000;
		8'h48		:	data	=	27'b001101001011111010000010000; //ADD ACC A
		8'h49		:	data	=	27'b000000000000000000000000000;
		8'h4A		:	data	=	27'b000000000000000000000000000;
		8'h4B		:	data	=	27'b000000000000000000000000000;
		8'h4C		:	data	=	27'b000000000000000000000000000;
		8'h4D		:	data	=	27'b000000000000000000000000000;
		8'h4E		:	data	=	27'b000000000000000000000000000;
		8'h4F		:	data	=	27'b000000000000000000000000000;
		8'h50		:	data	=	27'b000000000000000001000000000; //JMP CTE
		8'h51		:	data	=	27'b000000000000000000000100000;
		8'h52		:	data	=	27'b000000001000000010001010000;
		8'h53		:	data	=	27'b000000000000000000000000000;
		8'h54		:	data	=	27'b000000000000000000000000000;
		8'h55		:	data	=	27'b000000000000000000000000000;
		8'h56		:	data	=	27'b000000000000000000000000000;
		8'h57		:	data	=	27'b000000000000000000000000000;
		8'h58		:	data	=	27'b000000000000000001000000111; //JZ CTE
		8'h59		:	data	=	27'b000000000000000000000100000;
		8'h5A		:	data	=	27'b000000001000000010001010000;
		8'h5B		:	data	=	27'b000110001000000010000010000;
		8'h5C		:	data	=	27'b000000000000000000000000000;
		8'h5D		:	data	=	27'b000000000000000000000000000;
		8'h5E		:	data	=	27'b000000000000000000000000000;
		8'h5F		:	data	=	27'b000000000000000000000000000;
		8'h60		:	data	=	27'b000000000000000001000001011; //JN CTE
		8'h61		:	data	=	27'b000000000000000000000100000;
		8'h62		:	data	=	27'b000000001000000010001010000;
		8'h63		:	data	=	27'b000110001000000010000010000;
		8'h64		:	data	=	27'b000000000000000000000000000;
		8'h65		:	data	=	27'b000000000000000000000000000;
		8'h66		:	data	=	27'b000000000000000000000000000;
		8'h67		:	data	=	27'b000000000000000000000000000;
		8'h68		:	data	=	27'b000000000000000001000001111; //JC CTE
		8'h69		:	data	=	27'b000000000000000000000100000;
		8'h6A		:	data	=	27'b000000001000000010001010000;
		8'h6B		:	data	=	27'b000110001000000010000010000;
		8'h6C		:	data	=	27'b000000000000000000000000000;
		8'h6D		:	data	=	27'b000000000000000000000000000;
		8'h6E		:	data	=	27'b000000000000000000000000000;
		8'h6F		:	data	=	27'b000000000000000000000000000;
		8'h70		:	data	=	27'b000000000000000001000000000; //CALL DIR
		8'h71		:	data	=	27'b000110000000000000000100000;
		8'h72		:	data	=	27'b000000001000101000001000000;
		8'h73		:	data	=	27'b000000000001000001010000000;
		8'h74		:	data	=	27'b000000001101000000000000000;
		8'h75		:	data	=	27'b000111001001001000000000000;
		8'h76		:	data	=	27'b000110001001001000000000000;
		8'h77		:	data	=	27'b000111001001001010000010000;
		8'h78		:	data	=	27'b000110000001000001000000000; //RET
		8'h79		:	data	=	27'b000110001001001000000100000;
		8'h7A		:	data	=	27'b000000001000000010001010000;
		8'h7B		:	data	=	27'b000000000000000000000000000;
		8'h7C		:	data	=	27'b000000000000000000000000000;
		8'h7D		:	data	=	27'b000000000000000000000000000;
		8'h7E		:	data	=	27'b000000000000000000000000000;
		8'h7F		:	data	=	27'b000000000000000000000000000;
		8'h80		:	data	=	27'b000000000000000001000000000; //MOV ACC [DIR]
		8'h81		:	data	=	27'b000110001000000000000100000;
		8'h82		:	data	=	27'b000000000000000001001000000;
		8'h83		:	data	=	27'b000000000000000000000100000;
		8'h84		:	data	=	27'b000000001000111010001010000;
		8'h85		:	data	=	27'b000000000000000000000000000;
		8'h86		:	data	=	27'b000000000000000000000000000;
		8'h87		:	data	=	27'b000000000000000000000000000;
		8'h88		:	data	=	27'b000000000000000001000000000; //MOV DPTR CTE
		8'h89		:	data	=	27'b000110001000000000000100000;
		8'h8A		:	data	=	27'b000000001000010010001010000;
		8'h8B		:	data	=	27'b000000000000000000000000000;
		8'h8C		:	data	=	27'b000000000000000000000000000;
		8'h8D		:	data	=	27'b000000000000000000000000000;
		8'h8E		:	data	=	27'b000000000000000000000000000;
		8'h8F		:	data	=	27'b000000000000000000000000000;
		8'h90		:	data	=	27'b000000000000000001000000000; //AND ACC CTE
		8'h91		:	data	=	27'b000110001000000000000100000;
		8'h92		:	data	=	27'b000000001000101000001000000;
		8'h93		:	data	=	27'b001010001101111010000010000;
		8'h94		:	data	=	27'b000000000000000000000000000;
		8'h95		:	data	=	27'b000000000000000000000000000;
		8'h96		:	data	=	27'b000000000000000000000000000;
		8'h97		:	data	=	27'b000000000000000000000000000;
		8'h98		:	data	=	27'b001011001011111010000010000; //OR ACC A
		8'h99		:	data	=	27'b000000000000000000000000000;
		8'h9A		:	data	=	27'b000000000000000000000000000;
		8'h9B		:	data	=	27'b000000000000000000000000000;
		8'h9C		:	data	=	27'b000000000000000000000000000;
		8'h9D		:	data	=	27'b000000000000000000000000000;
		8'h9E		:	data	=	27'b000000000000000000000000000;
		8'h9F		:	data	=	27'b000000000000000000000000000;
		8'hA0		:	data	=	27'b001100001011111010000010000; //XOR ACC A
		8'hA1		:	data	=	27'b000000000000000000000000000;
		8'hA2		:	data	=	27'b000000000000000000000000000;
		8'hA3		:	data	=	27'b000000000000000000000000000;
		8'hA4		:	data	=	27'b000000000000000000000000000;
		8'hA5		:	data	=	27'b000000000000000000000000000;
		8'hA6		:	data	=	27'b000000000000000000000000000;
		8'hA7		:	data	=	27'b000000000000000000000000000;
		8'hA8		:	data	=	27'b001111001111111010000010000; //CA2 ACC
		8'hA9		:	data	=	27'b000000000000000000000000000;
		8'hAA		:	data	=	27'b000000000000000000000000000;
		8'hAB		:	data	=	27'b000000000000000000000000000;
		8'hAC		:	data	=	27'b000000000000000000000000000;
		8'hAD		:	data	=	27'b000000000000000000000000000;
		8'hAE		:	data	=	27'b000000000000000000000000000;
		8'hAF		:	data	=	27'b000000000000000000000000000;
		8'hB0		:	data	=	27'b001111001011011010000010000; //CA2 A
		8'hB1		:	data	=	27'b000000000000000000000000000;
		8'hB2		:	data	=	27'b000000000000000000000000000;
		8'hB3		:	data	=	27'b000000000000000000000000000;
		8'hB4		:	data	=	27'b000000000000000000000000000;
		8'hB5		:	data	=	27'b000000000000000000000000000;
		8'hB6		:	data	=	27'b000000000000000000000000000;
		8'hB7		:	data	=	27'b000000000000000000000000000;
		8'hB8		:	data	=	27'b001000011111111010000010000; //SLR ACC
		8'hB9		:	data	=	27'b000000000000000000000000000;
		8'hBA		:	data	=	27'b000000000000000000000000000;
		8'hBB		:	data	=	27'b000000000000000000000000000;
		8'hBC		:	data	=	27'b000000000000000000000000000;
		8'hBD		:	data	=	27'b000000000000000000000000000;
		8'hBE		:	data	=	27'b000000000000000000000000000;
		8'hBF		:	data	=	27'b000000000000000000000000000;
		8'hC0		:	data	=	27'b001000101111111010000010000; //SLL ACC
		8'hC1		:	data	=	27'b000000000000000000000000000;
		8'hC2		:	data	=	27'b000000000000000000000000000;
		8'hC3		:	data	=	27'b000000000000000000000000000;
		8'hC4		:	data	=	27'b000000000000000000000000000;
		8'hC5		:	data	=	27'b000000000000000000000000000;
		8'hC6		:	data	=	27'b000000000000000000000000000;
		8'hC7		:	data	=	27'b000000000000000000000000000;
		8'hC8		:	data	=	27'b001110001111111010000010000; //INC ACC
		8'hC9		:	data	=	27'b000000000000000000000000000;
		8'hCA		:	data	=	27'b000000000000000000000000000;
		8'hCB		:	data	=	27'b000000000000000000000000000;
		8'hCC		:	data	=	27'b000000000000000000000000000;
		8'hCD		:	data	=	27'b000000000000000000000000000;
		8'hCE		:	data	=	27'b000000000000000000000000000;
		8'hCF		:	data	=	27'b000000000000000000000000000;
		8'hD0		:	data	=	27'b000000000000000000000000000; // MOV [DIR] ACC
		8'hD1		:	data	=	27'b000000000000000000000000000;
		8'hD2		:	data	=	27'b000000000000000000000000000;
		8'hD3		:	data	=	27'b000000000000000000000000000;
		8'hD4		:	data	=	27'b000000000000000000000000000;
		8'hD5		:	data	=	27'b000000000000000000000000000;
		8'hD6		:	data	=	27'b000000000000000000000000000;
		8'hD7		:	data	=	27'b000000000000000000000000000;
		8'hD8		:	data	=	27'b000000000000000000000000000; //
		8'hD9		:	data	=	27'b000000000000000000000000000;
		8'hDA		:	data	=	27'b000000000000000000000000000;
		8'hDB		:	data	=	27'b000000000000000000000000000;
		8'hDC		:	data	=	27'b000000000000000000000000000;
		8'hDD		:	data	=	27'b000000000000000000000000000;
		8'hDE		:	data	=	27'b000000000000000000000000000;
		8'hDF		:	data	=	27'b000000000000000000000000000;
		8'hE0		:	data	=	27'b000000000000000000000000000; //
		8'hE1		:	data	=	27'b000000000000000000000000000;
		8'hE2		:	data	=	27'b000000000000000000000000000;
		8'hE3		:	data	=	27'b000000000000000000000000000;
		8'hE4		:	data	=	27'b000000000000000000000000000;
		8'hE5		:	data	=	27'b000000000000000000000000000;
		8'hE6		:	data	=	27'b000000000000000000000000000;
		8'hE7		:	data	=	27'b000000000000000000000000000;
		8'hE8		:	data	=	27'b000000000000000000000000000; //
		8'hE9		:	data	=	27'b000000000000000000000000000;
		8'hEA		:	data	=	27'b000000000000000000000000000;
		8'hEB		:	data	=	27'b000000000000000000000000000;
		8'hEC		:	data	=	27'b000000000000000000000000000;
		8'hED		:	data	=	27'b000000000000000000000000000;
		8'hEE		:	data	=	27'b000000000000000000000000000;
		8'hEF		:	data	=	27'b000000000000000000000000000;
		8'hF0		:	data	=	27'b000000000000000000000000000; //
		8'hF1		:	data	=	27'b000000000000000000000000000;
		8'hF2		:	data	=	27'b000000000000000000000000000;
		8'hF3		:	data	=	27'b000000000000000000000000000;
		8'hF4		:	data	=	27'b000000000000000000000000000;
		8'hF5		:	data	=	27'b000000000000000000000000000;
		8'hF6		:	data	=	27'b000000000000000000000000000;
		8'hF7		:	data	=	27'b000000000000000000000000000;
		8'hF8		:	data	=	27'b000000000000000000000000000; //
		8'hF9		:	data	=	27'b000000000000000000000000000;
		8'hFA		:	data	=	27'b000000000000000000000000000;
		8'hFB		:	data	=	27'b000000000000000000000000000;
		8'hFC		:	data	=	27'b000000000000000000000000000;
		8'hFD		:	data	=	27'b000000000000000000000000000;
		8'hFE		:	data	=	27'b000000000000000000000000000;
		8'hFF		:	data	=	27'b000000000000000000000000000;
		default	:	data	=	27'b000000000000000000000000000;
	endcase

endmodule